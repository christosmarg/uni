library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity instrmem is port (
	addr:	in std_logic_vector(31 downto 0);
	c:	out std_logic_vector(31 downto 0)
);
end instrmem;

architecture dataflow of instrmem is

type instr_arr is array(0 to 31) of std_logic_vector (31 downto 0);
constant instr_mem: instr_arr := (
	"00000000010001100010000000100000", -- 0 add $4, $2, $6
	"00000000010001100010100000100010", -- 1 sub $5, $2, $6
	"11111100100001010000000000000000", -- 2 read $4, $5
	"00000000000000000000000000000000", -- 3
	"00000000000000000000000000000000", -- 4
	"00000000000000000000000000000000", -- 5
	"00000000000000000000000000000000", -- 6
	"00000000000000000000000000000000", -- 7
	"00000000000000000000000000000000", -- 8
	"00000000000000000000000000000000", -- 9
	"00000000000000000000000000000000", -- 10
	"00000000000000000000000000000000", -- 11
	"00000000000000000000000000000000", -- 12
	"00000000000000000000000000000000", -- 13
	"00000000000000000000000000000000", -- 14
	"00000000000000000000000000000000", -- 15
	"00000000000000000000000000000000", -- 16
	"00000000000000000000000000000000", -- 17
	"00000000000000000000000000000000", -- 18
	"00000000000000000000000000000000", -- 19
	"00000000000000000000000000000000", -- 20
	"00000000000000000000000000000000", -- 21
	"00000000000000000000000000000000", -- 22
	"00000000000000000000000000000000", -- 23
	"00000000000000000000000000000000", -- 24
	"00000000000000000000000000000000", -- 25
	"00000000000000000000000000000000", -- 26
	"00000000000000000000000000000000", -- 27
	"00000000000000000000000000000000", -- 28
	"00000000000000000000000000000000", -- 29
	"00000000000000000000000000000000", -- 30
	"00000000000000000000000000000000"  -- 31
);

begin
	-- Our addresses are multiples of 4, so ignore the last 2 bits.
	c <= instr_mem(to_integer(unsigned(addr(31 downto 2))));
end dataflow;
