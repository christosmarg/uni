library ieee;
use ieee.std_logic_1164.all;

entity pc is port (
);
end pc;

architecture behav of pc is
begin
end behav;
