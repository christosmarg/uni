library ieee;
use ieee.std_logic_1164.all;

entity adder32 is port (
);
end adder32;

architecture behav of adder32 is

begin
end behav;
