library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity instrmem is port (
	addr:	in std_logic_vector(3 downto 0);
	c:	out std_logic_vector(31 downto 0)
);
end instrmem;

architecture dataflow of instrmem is

type instr_arr is array(0 to 15) of std_logic_vector (31 downto 0);
constant instr_mem: instr_arr := (
	"11111111111111111111111111111111", -- 0
	"10001010100101010101000011101111", -- 1
	"11111111111111111111111111111111", -- 2
	"00000000000000000000000000000000", -- 3
	"11111111111111111111111111111111", -- 4
	"00000000000000000000000000000000", -- 5
	"00000000101001100010000000100000", -- 6
	"11111111111111111111111111111111", -- 7
	"11111111111111111111111111111111", -- 8
	"11111111111111111111111111111111", -- 9
	"10101010101011110000101110001010", -- 10
	"11111111111111100000000000000000", -- 11
	"10001011101010111010111101010111", -- 12
	"11111111111111111111111111111111", -- 13
	"10110111000111010101010101111111", -- 14
	"11111111111111111111111111111111"  -- 15
);

begin
	c <= instr_mem(to_integer(unsigned(addr)));
end dataflow;
