library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity instrmem is port (
	addr:	in std_logic_vector(3 downto 0);
	c:	out std_logic_vector(31 downto 0)
);
end instrmem;

architecture dataflow of instrmem is

type instr_arr is array(0 to 15) of std_logic_vector (31 downto 0);
constant instr_mem: instr_arr := (
	"00000000000000000000000000000000", -- 0
	"00000000000000000000000000000000", -- 1
	"00000000000000000000000000000000", -- 2
	"00000000000000000000000000000000", -- 3
	"00000000000000000000000000000000", -- 4
	"00000000000000000000000000000000", -- 5
	"00000000000000000000000000000000", -- 6
	"00000000000000000000000000000000", -- 7
	"00000000000000000000000000000000", -- 8
	"00000000000000000000000000000000", -- 9
	"00000000000000000000000000000000", -- 10
	"00000000000000000000000000000000", -- 11
	"00000000000000000000000000000000", -- 12
	"00000000000000000000000000000000", -- 13
	"00000000000000000000000000000000", -- 14
	"00000000000000000000000000000000"  -- 15
);

begin
	c <= instr_mem(to_integer(unsigned(addr)));
end dataflow;
